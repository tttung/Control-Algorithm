`timescale 1ns / 1ps
/**********************************************************************************
;** ��������: filter.v
;** ��������: ȥ���ź���ë�̣�С��2��ʱ��cp������źţ�
;** �䡡��:   cp    :ʱ���ź�
;**           x_in  :����ë�̵��ź�
;** �䡡�� :  y_out :ȥ��ë�̺���ź�
;** ȫ�ֱ���: y_out
;** ����ģ��: ��
;**-------------------------------------------------------------------------------*/

module filter ( cp, x_in,y_out);
  // �˿�����
     input cp;                   // ����ʱ�����   
     input x_in;                 // ����ǰ�����ź�
     output y_out;               // ����������ź�

  // �˿ڱ������Ͷ���
     wire cp;                    // ������Ϊinput��inout�͵ı���ֻ�ܱ�����Ϊ������
     wire x_in;                  // �����ͱ����������ӹ�ϵ
     reg y_out;                  // y_outΪ����Ĵ�������
  
  // �ڲ��Ĵ�������
     reg [1:0] q;                // ����һ��1λ��3��Ԫ�ص����黺��Ĵ���
     reg [1:0] sum;              // ������ͼĴ���
     integer i;                  // ��������

  // ��������
     always @(posedge cp)        // ������ô������ݻ�����
          begin
          //     q[2] = q[1];
               q[1] = q[0];
               q[0] = x_in;
          end
     always @(posedge cp)
          begin
               sum = 0;
               for(i=0;i<2;i=i+1)
               begin
                   if (q[i] == 1)
                       sum = sum +1;
                   else
                       sum = sum;
               end
               if (sum > 1)     // ����1��ʱ��������ź���Ϊ����ë���ź�
                   y_out <= 1;
               else
                   y_out <= 0;
           end 

  endmodule


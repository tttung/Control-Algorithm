`timescale 1ns / 1ps
/**--------------�ļ���Ϣ------------------------------------------------------------------------------
;**��   ��   ��: pwm.v
;**��        ��: Verilog HDL������EPM7128STC100-10�ϣ�������·����180����λ��PWM�źš���PWM�źž���
;**              ��ë�̴����ڹ�������ѹ�͹��ȱ���ʱ���Զ��ر�PWM�źš���MAX+plusII10.1���롣
;**--------------��ʷ�汾��Ϣ--------------------------------------------------------------------------
;** ��  ��: V1.1
;**         ����V1.0ռ�õ��߼���̫��ֻ����2500��оƬ��ʵ�֣��ʸı�PWM�㷨������1200��оƬ��ʵ��
;**--------------��ʷ�汾��Ϣ--------------------------------------------------------------------------
;** ��  ��: V1.2
;**         ��������ʱ,PWM-A,PWM-B��ͬ������ռ�ձ�1300��
;**---------------------------------------------------------------------------------------------------*/

module pwm (clock,data_in,pwm_out,rst_n);
  // �˿�����
     input clock;                          // ����ʱ����˿�
	  input rst_n;
     input[11:0] data_in;                   // ����12λ����������˿�
     output pwm_out;                     // ����PWM_A����˿�

  // �˿ڱ������Ͷ���
                               // ������Ϊinput��inout�͵ı���ֻ�ܱ�����Ϊ������
     wire[11:0] data_in;                                    
     wire  pwm_out;                       // PWM_A����Ĵ�������
	 
	 // wire clock; 
                                           // ��output�Ͷ˿�������Ӷ�����Ĭ��Ϊwire��
	  
  // �ڲ��Ĵ�������
     reg[12:0] counter1;                    // ʱ�Ӽ����Ĵ���,��ʼֵĬ����0 
  //   reg[11:0] counter2;  
  //   reg flag ;                            // ��־�Ĵ���,��ʼֵĬ����0 
     reg pwm_A;

  // ��������
     always @(posedge clock)               
                                           // ����clock�ź������ش���
                                           // (2500*2)*40KHz=200MHz��clock�źţ�����160KHz���ǲ�
        // begin
             
          //   if (flag == 1)                // ����������ǲ�����б��
         //    begin 
          //        if (counter2 < 2500)
          //            counter2 <= counter2 + 1;
          //        else
          //       begin
          //             counter2 <= 0;
          //             flag <= 0;          // ��ǰ���������ǲ�����б�±�־
          //        end
          //   end
          //   else                          // ǰ���������ǲ�����б��
             begin
                  if (counter1 < 5000)      // ��������Ϊ5.4us
                      counter1 <= counter1 + 1;                  
                  else     
                  begin
                       counter1 <= 0;
                     //  flag <= 1;          // �����������ǲ�����б�±�־
                  end

             end 
       //  end

     always @(counter1) // or counter2
        // begin
           //  begin
             //     if(flag==0)
                  begin
                       if(counter1 < 3500)
                            pwm_A <= 1;        // �ǣ�������ߵ�ƽ
                       else
                            pwm_A <= 0;        // ��������͵�ƽ
                  end
						//else
                 // begin
                 //      if(counter2 < 150)
                  //          pwm_A <= 1;        // �ǣ�������ߵ�ƽ
                  //     else
                  //          pwm_A <= 0;        // ��������͵�ƽ
                //  end
          //   end
        // end
         
     filter U1(.cp(clock),.x_in(pwm_A),.y_out(pwm_out)); // ����PWM-A�˲�ģ�� 
 
 endmodule


